module test_fifo #(
) (
);
  logic [ 7:0] rx_buf[ 7:0];
  logic [ 4:0] rx_rptr;
  logic [ 4:0] rx_wptr;
endmodule